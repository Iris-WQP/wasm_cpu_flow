`define log2_S 5
`define log2_Width_max 10
`define log2_Height_max 10

`define MAX_DW    8                 // datawidth
`define MAX_log2DW   3

`define MAX_DW2 (`MAX_DW*2)

`define Tin 8
`define log2_Tin 3

`define Tout 8
`define log2_Tout 3

`define Acc_Delay 4
`define Acc_Height_Num 256
`define Tin_Acc_Delay `log2_Tin